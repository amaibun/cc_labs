library verilog;
use verilog.vl_types.all;
entity tb_demux1to8 is
end tb_demux1to8;
